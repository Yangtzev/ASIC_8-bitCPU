`timescale 1 ns / 1ns
module mem ( data, addr, read, write );
input [7:0] data;
input [7:0] addr;
input read;
input write;

reg [7:0] memory [0:31];

assign data= (read)?memory[addr]:8'hZ;

always @(posedge write)
begin
memory[addr]<=data[7:0];
end

endmodule
